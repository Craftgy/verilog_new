module async_fifo #(
    parameter DATA_WIDTH = 4;
    p
);

endmodule