module sync_fifo # (
    parameter DATA_WIDTH = 8,
    p
);
    
endmodule