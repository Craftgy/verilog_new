module SPI #(
    parameter CMD_WIDTH,
    par
) (
    ports
);
    
endmodule