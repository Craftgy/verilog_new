module sync_fifo # (
     DATA_WIDTH = 8,
    parameter
);
    
endmodule