module sync_fifo # (
    par
);
    
endmodule