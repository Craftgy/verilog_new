module s();

endmodule