module CRCCYC