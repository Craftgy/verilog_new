module CRCCYC(Clock,Data_)