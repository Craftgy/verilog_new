module sysnv();

endmodule