module SPI #(
    parameter W
) (
    ports
);
    
endmodule