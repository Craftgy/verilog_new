module Redge(
    clk,
    din,
    pulse
);
input clk