module sync_fifo # (
    ports
);
    
endmodule