module sync_fifo # (
    parameter DATA_W
);
    
endmodule