module async();

endmodule