module sync_fifo # (
    
);
    
endmodule