module Redge(
    clk,
    din,
    pulse
);