module async_fifo #(
    parameter DATA_WIDTH = 4;
    parameter FIFO_DEPTH = 16;
);

endmodule