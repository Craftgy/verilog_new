module Redge(
    clk,
    
)