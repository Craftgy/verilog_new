module Redge(
    clk,
    din,
    
)