module sync_fio (
    ports
);
    
endmodule