module SPI #(
    parameter CMD_W
) (
    ports
);
    
endmodule