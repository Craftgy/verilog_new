module Redge(
    
)