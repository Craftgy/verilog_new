module SPI #(
    parameter CMD_WIDTH,
) (
    ports
);
    
endmodule