module sync_fi (
    ports
);
    
endmodule