module Redge(
    clk,
)