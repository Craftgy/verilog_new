module CRCC