module async_fifo #(
    par
);

endmodule