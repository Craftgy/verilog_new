module CRCCYC(Clock,)