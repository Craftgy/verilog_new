module R