module Redge(
    clk,
    din
)