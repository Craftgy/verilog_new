module CRCCYC()