module sync_F (
    ports
);
    
endmodule