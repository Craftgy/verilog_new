module sysc();

endmodule