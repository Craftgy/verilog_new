module SPI #(
    parameter CMD_WIDTH = 12,
    parameter  = 
) (
    ports
);
    
endmodule