module CRCCYC(Clock,Data_IN,CRC_En)