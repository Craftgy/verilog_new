module sysn();

endmodule