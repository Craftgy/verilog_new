module async_fifo #(
    parameter DATA_WIDTH = ;
);

endmodule