module Redge()