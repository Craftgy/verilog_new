module Redge(
    clk,
    din,
    pulse
);
input wire clk