module CRCCYC(Clock,Data_IN,CRC_En,CRC_Clr,CRC_Out);
input 