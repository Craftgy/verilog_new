module SPI #(
    parameters
) (
    ports
);
    
endmodule