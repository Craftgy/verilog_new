module Redge(
    clk,
    din,
    pu
)