module Redge(
    in
)