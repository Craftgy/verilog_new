module CRCCYC(Clock,Data_IN)