module SPI #(
    parameter CMD_WIDTH = ,
    parameter  = 
) (
    ports
);
    
endmodule