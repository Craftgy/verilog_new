module sysc_fifo_tb();

endmodule