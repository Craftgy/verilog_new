module async_fifo #();

endmodule