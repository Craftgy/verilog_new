module async_fifo #(
    parameter DATA = ;
);

endmodule