module Redge