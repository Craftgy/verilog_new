module SPI #(
    parameter CMD_WIDTH,
    pa
) (
    ports
);
    
endmodule