module async_fifo #(
    parameter  = ;
);

endmodule