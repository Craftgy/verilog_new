module SPI #(
    parameter CMD_WIDTH = 12,
    parameter READ_WIDTH = 
) (
    ports
);
    
endmodule