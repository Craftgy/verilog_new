module SPI #(
    parameter 
) (
    ports
);
    
endmodule