module SPI #(
    parameter CMD_WIDTH = 12,
    parameter READ_WIDTH = 8,
) (
    ports
);
    
endmodule