module sync_fifo # (
    parameter DATA
);
    
endmodule