module CRCCYC(Clock,Data)