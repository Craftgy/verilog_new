module Redge(
    clk
)