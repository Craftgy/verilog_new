module sync (
    ports
);
    
endmodule